interface and_intf();
bit a;
bit b;
bit y;

endinterface
