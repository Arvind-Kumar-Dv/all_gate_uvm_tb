typedef uvm_sequencer#(and_tx) and_sqr;
